library verilog;
use verilog.vl_types.all;
entity CONTROL_UNITY_vlg_vec_tst is
end CONTROL_UNITY_vlg_vec_tst;
