library verilog;
use verilog.vl_types.all;
entity SHIFTER_vlg_vec_tst is
end SHIFTER_vlg_vec_tst;
